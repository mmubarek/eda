package RISC_ISA_pkg;
  parameter INSTR_WIDTH = 32;
  parameter DATA_WIDTH = 32;
  parameter ADDR_WIDTH = 32;
  parameter REG_ADDR_WIDTH = 5;
  parameter REG_COUNT = 32;
  localparam OP_R_TYPE = 7'b0110011;
  localparam OP_I_TYPE_ARITH = 7'b0010011;
  localparam OP_LOAD = 7'b0000011;
  localparam OP_STORE = 7'b0100011;
  localparam OP_BRANCH = 7'b1100011;
  localparam FUNCT3_ADD_SUB_ADDI = 3'b000;
  localparam FUNCT3_LW_SW = 3'b010;
  localparam FUNCT3_BEQ = 3'b000;
  localparam FUNCT7_ADD = 7'b0000000;
  localparam FUNCT7_SUB = 7'b0100000;
  localparam ALU_ADD = 3'b000;
  localparam ALU_SUB = 3'b001;
  localparam ALU_PASS_B = 3'b010;
  localparam ALU_EQ_CHECK = 3'b011;
  localparam PC_SRC_INC = 2'b00;
  localparam PC_SRC_BRANCH = 2'b01;
  localparam ALU_SRC_A_REG = 1'b0;
  localparam ALU_SRC_A_PC = 1'b1;
  localparam ALU_SRC_B_REG = 1'b0;
  localparam ALU_SRC_B_IMM = 1'b1;
  localparam IMM_TYPE_I = 2'b00;
  localparam IMM_TYPE_S = 2'b01;
  localparam IMM_TYPE_B = 2'b10;
  localparam WB_SRC_ALU = 2'b00;
  localparam WB_SRC_MEM = 2'b01;
endpackage